`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:47:58 06/08/2019 
// Design Name: 
// Module Name:    rom_data1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module rom_data1(
    adder_1    ,
    
    //�����ź�,����dout
    data_1    );

    //��������
    

    //�����źŶ���
    input [5:0]          adder_1  ;
  

    //����źŶ���
    output[507:0]         data_1   ;

    //����ź�reg����
    reg   [507:0]         data_1   ;

   

    //����߼�д��
    always@(*)begin 
        case(adder_1)
			 6'd1 :    data_1 = 508'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
 6'd2 :    data_1 = 508'h000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000003000000000000;
 6'd3 :    data_1 = 508'h000000FC00000001F00000000000200000000000000003000000001F0001FA000000000000000000000003C000000000000000000F00000003FE0000000000;
 6'd4 :    data_1 = 508'h000001FF00000301FE00000000001F000000000000000FE00000001FE001FC000000000380000000000000FE00000000000000000FF8000003F80000000000;
 6'd5 :    data_1 = 508'h000001F800001FC1F000000000001FFFFFFFFFFFFFFFFFF00000001F8001F8000000007FE00000000000003FC0000000000000000FC0000003F00000000000;
 6'd6 :    data_1 = 508'h000003F00001FFF1F03E000000001F00007C0001F0000FC00000001F8001F8000C003FFFF80000000000001FE0000000000000000F80000003F00000000000;
 6'd7 :    data_1 = 508'h000007E0001FF801F007E00000001F00007C0001F0000FC00000000F8001F8000FFFE0000000000000000007E0000000000000000F80000003F00000000000;
 6'd8 :    data_1 = 508'h00000F8003FF8001F001FC0000001F00007C0001F0000FC00000000F8001F8780F8000000000000000000003C0000000180000000F80000003F00000000000;
 6'd9 :    data_1 = 508'h00001F01FC0F8001F0007E0000001F00007C0001F0000FC00001FFFFFFFFFFFF0F800000000000000000000100000000FE0000000F80000003F00000000000;
 6'd10 :    data_1 = 508'h00003E00000F8001F0003E0000001F00007C0001F0000FC00000000F8001F8000F8000000000FFFFFFFFFFFFFFFFFFFFFFC000000F80000003F00007C00000;
 6'd11 :    data_1 = 508'h00007C00000F8001F000180000001F00007C0001F0000FC00000000F8001F8000F80000000001F80000003F000000000002000000F8003FFFFFFFFFFF80000;
 6'd12 :    data_1 = 508'h0000FC00000F8001F800000000001F00007C0001F0000FC00000000F8001F8000F80000000000000000003F000000000000000000F8000C003F00007E00000;
 6'd13 :    data_1 = 508'h0001FF80000F8000F8000F8000001F00007C0001F0000FC00000000F8001F8000F80000000000000000003F000000000000000000F807C0003F00007C00000;
 6'd14 :    data_1 = 508'h0003FE10000F8000F8003FF000001FFFFFFFFFFFFFFFFFC00000000FFFFFF8000F80000000000000000003E00000000000000FFFFFFFFF8003F00007C00000;
 6'd15 :    data_1 = 508'h0007BE0FFFFFFFFFFFFFC00800001F000003E00000000FC00000000F8001F8000F80000040000000000007E000000000000001E00F80004003F00007C00000;
 6'd16 :    data_1 = 508'h001F3E00000F8000F800000000001F00000FFE00000008000000000F8001F8000F800003F0000000000007E000000000000000000F80000003F00007C00000;
 6'd17 :    data_1 = 508'h003C3E00000F8000F800180000002000003FE000000000000000000F8001F8000FFFFFFFFE000000000007C000000780000000000F80000003F00007C00000;
 6'd18 :    data_1 = 508'h00703E00000F8000F8003F8000000000007F0000000700000000000F8001F8000F8001F00000000000000FFFFFFFFFF8000000000F80000003E00007C00000;
 6'd19 :    data_1 = 508'h01C03E00000F8000F8007FC00000000001FC0000001FE0000000000F8001F8000F8001F00000000000000FC000000FF0000000000F80000003E00007C00000;
 6'd20 :    data_1 = 508'h03003E00000F80F0F800FE000000000007F3FFFFFFFFF8000000000FFFFFF8000F8001F00000000000001F8000001FC0000000000F80000003E00007C00000;
 6'd21 :    data_1 = 508'h0C003E00000F9F007C01F800000000003F800000003F80000000000F8001F8000F8001F00000000000001F0000001F80000000000F80000003E00007C3E000;
 6'd22 :    data_1 = 508'h00003E00000FF8007C03F00000000000FC00000000FE00000000000F8001F8000F8001F00000000000003F0000001F80000000000F83FFFFFFFFFFFFFFFC00;
 6'd23 :    data_1 = 508'h00003E0000FF80007E07C00000000007FF00000001FC00000000000F8001F8000F8001F00000000000007E0000001F80000000000F807E0007E60000000200;
 6'd24 :    data_1 = 508'h00003E001FFF80003E1F80000000003F83F0000007F000000000000F8001F8781F8001F0000000000000FC0000003F00000000000F80000007C30000000000;
 6'd25 :    data_1 = 508'h00003E0FFF0F80003F3E0000000001F800FE00001FC00000000FFFFFFFFFFFFE1F8001F0000000000001F80000003F00000000000F8000000FC18000000000;
 6'd26 :    data_1 = 508'h00003E0FF00F80001FFC000000000F80007F80007F0000000001C000000000011F0001F0000000000003F00000003F00000000000F8000001F81E000000000;
 6'd27 :    data_1 = 508'h00003E03800F80000FF000000000F000001F8001FC00000000000000000000003F0001F0000000000007C00000007E00000000000F80FFC01F00F000000000;
 6'd28 :    data_1 = 508'h00003E00000F800007C00018000F0000000F800FF000000000000001800E00003E0001F000000000001F800000007E00000000000FFF80007E007C00000000;
 6'd29 :    data_1 = 508'h00003E00000F80001FF0003000000000000F007F8000000000000003F003F0007C0001F000000000003E00000000FC000000003FFFE00000FC001E00000000;
 6'd30 :    data_1 = 508'h00003E00000F8000FDF8007000000000000003FC0000000000000007F800FE00F80001F00000000000F800000000FC00000007FFF0000001F8000F80000000;
 6'd31 :    data_1 = 508'h00003E00000F8003E07E00F00000000000001FE0000000000000001FC0003F01F00001F00000000003E000000001FC00000003FC00000007E00003F0000000;
 6'd32 :    data_1 = 508'h00003E00000F801F003F80F0000000000003FE00000000000000003E00001F83E00001F0000000000F8000000001F800000000C00000001F800001FC000000;
 6'd33 :    data_1 = 508'h00003E00000F8070000FF1E000000000003FE00000000000000000F800000F0F800001F0000000003E0000000003F80000000000000000FC0000007FC00000;
 6'd34 :    data_1 = 508'h00003E03801F83800003FFE0000000000FFC000000000000000003E00000061E000001F000000001F000003F0007F00000000000000007E00000001FFC0000;
 6'd35 :    data_1 = 508'h00003E007FFF800000007FF000000003FE0000000000000000000F0000000078000001F00000000F80000001FFFFE0000000000000007E0000000003FFF000;
 6'd36 :    data_1 = 508'h00003E0003FE000000000FF0000003FE000000000000000000007800000001C0000001F000000078000000003FFF8000000000000007E00000000000FFFF00;
 6'd37 :    data_1 = 508'h00003E0000F8000000000070003FFC0000000000000000000001C00000000E00000001F000000F800000000007FC00000000000000FC0000000000001F8000;
 6'd38 :    data_1 = 508'h000030000000000000000000000000000000000000000000000000000000300000000180000010000000000003000000000000000F00000000000000020000;
 6'd39 :    data_1 = 508'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
 6'd40 :    data_1 = 508'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
							

default:   data_1 = 508'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

      endcase
    
   end
   endmodule
